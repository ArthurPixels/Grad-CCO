library ieee;
use ieee.std_logic_1164.all;

entity map3 is
	port
	(
		F0, F1, F2, F3, F4, F5, F6, F7, F8, F9, F10, F11, F12, F13, F14, F15: out std_logic_vector(31 downto 0)
	);
end map3;	
	
architecture map3_struct of map3 is
begin
	F0  <= "00000000000000000000000000000000";
	F1  <= "00000000000000000000000000000000";
	F2  <= "00000000000000000000000000000000";
	F3  <= "00000000111100000001111000000000";
	F4  <= "00000000100100000001001000000000";
	F5  <= "00000000111100000001111000000000";
	F6  <= "00000000000000000000000000000000";
	F7  <= "00000000010000000000010000000000";
	F8  <= "00000000010000000000010000000000";
	F9  <= "00000000001000000000100000000000";
	F10 <= "00000000000111111110000000000000";
	F11 <= "00000000000000000000000000000000";
	F12 <= "00000000000000000000000000000000";
	F13 <= "00000000000000000000000000000000";
	F14 <= "00000000000000000000000000000000";
	F15 <= "00000000000000000000000000000000";
end map3_struct;