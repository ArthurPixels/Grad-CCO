library ieee;
use ieee.std_logic_1164.all;

entity map4 is
	port
	(
		F0, F1, F2, F3, F4, F5, F6, F7, F8, F9, F10, F11, F12, F13, F14, F15: out std_logic_vector(31 downto 0)
	);
end map4;	
	
architecture map4_struct of map4 is
begin
	F0  <= "00000111100110001001110000000000";
	F1  <= "00000100000101001001001000000000";
	F2  <= "00000111111100111101000100000000";
	F3  <= "00000000000100011001001000000000";
	F4  <= "00000000000100001111110000000000";
	F5  <= "00000001000000000000000000000000";
	F6  <= "00000000000000000000010000000000";
	F7  <= "11111100000000000000000000000000";
	F8  <= "10100100100000000000000000000000";
	F9  <= "11111111111111111000001111111111";
	F10 <= "10000000000001000000000000000000";
	F11 <= "11111100011110000000000111001011";
	F12 <= "00000000000000000000000000010000";
	F13 <= "00000000000000000000000000010000";
	F14 <= "00000000000000000000000000010000";
	F15 <= "00000000000000000000000000010000";
end map4_struct;